//*****************************************************************************
// qwic51_defs.vh
//
// This module is the global defines of qwic51.
//
// Change History:
//  VER.   Author         DATE              Change Description
//  0.1    Qiwei Wu       Nov. 24, 2019     Initial Release
//
//*****************************************************************************
// Define
`define CPU_DATA_WIDTH 8
`define CPU_ADDR_WIDTH 8
`define CPU_RAM_ADDWID 8
`define CPU_ROM_ADDWID 8
