//*****************************************************************************
// qwic51_include.vh
//
// This module is the includes defines of qwic51.
//
// Change History:
//  VER.   Author         DATE              Change Description
//  0.1    Qiwei Wu       Nov. 30, 2019     Initial Release
//
//*****************************************************************************

`include "qwic51_defs.vh"
`include "qwic51_memdefs.vh"
`include "qwic51_arithmeticdefs.vh"
`include "qwic51_instructdefs.vh"